string s1 = "Hello World";

$display("%s", s1);
